
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;

entity Register_Banc is
    Port ( ADD : in  STD_LOGIC_VECTOR (7 downto 0);
			  IND : in STD_LOGIC_VECTOR (2 downto 0);
           DAT : in  STD_LOGIC_VECTOR (7 downto 0);
           RX_E : in  STD_LOGIC;
           TX_E : in  STD_LOGIC;
			  Reset : in STD_LOGIC;
           D_TX : out  STD_LOGIC);
end Register_Banc;

architecture Behavioral of Register_Banc is
type memoire is array (0 to 255) of STD_LOGIC_VECTOR (7 downto 0);
	signal registery : memoire := 
		(X"AA",X"44",X"33",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00") ;
	
begin

process(ADD,RX_E,Reset)
begin
	if Reset='1' and Reset'event
	then
		for i in 0 to 255  loop
			registery(i)<= X"00" ;
		end loop  ;
	end if;
	if RX_E='1' and Reset='0'
	then
		registery(conv_integer(ADD)) <= DAT ;
	end if;
end process;

process(ADD,IND,TX_E,Reset)
begin
	if TX_E='1' and Reset='0'
	then
		D_TX <= registery(conv_integer(ADD))(conv_integer(IND)) ;
	end if;
end process;

end Behavioral;

